library verilog;
use verilog.vl_types.all;
entity ProgramCounter_vlg_vec_tst is
end ProgramCounter_vlg_vec_tst;
