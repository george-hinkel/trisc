library verilog;
use verilog.vl_types.all;
entity PartBController_vlg_vec_tst is
end PartBController_vlg_vec_tst;
