library verilog;
use verilog.vl_types.all;
entity Lab1_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab1_vlg_check_tst;
