library verilog;
use verilog.vl_types.all;
entity RippleCarryAdder_vlg_vec_tst is
end RippleCarryAdder_vlg_vec_tst;
